module Systolic_Array10x10 (
	output reg [31:0]
		 out0_0, out0_1, out0_2, out0_3, out0_4, out0_5, out0_6, out0_7, out0_8, out0_9,
		 out1_0, out1_1, out1_2, out1_3, out1_4, out1_5, out1_6, out1_7, out1_8, out1_9,
		 out2_0, out2_1, out2_2, out2_3, out2_4, out2_5, out2_6, out2_7, out2_8, out2_9,
		 out3_0, out3_1, out3_2, out3_3, out3_4, out3_5, out3_6, out3_7, out3_8, out3_9,
		 out4_0, out4_1, out4_2, out4_3, out4_4, out4_5, out4_6, out4_7, out4_8, out4_9,
		 out5_0, out5_1, out5_2, out5_3, out5_4, out5_5, out5_6, out5_7, out5_8, out5_9,
		 out6_0, out6_1, out6_2, out6_3, out6_4, out6_5, out6_6, out6_7, out6_8, out6_9,
		 out7_0, out7_1, out7_2, out7_3, out7_4, out7_5, out7_6, out7_7, out7_8, out7_9,
		 out8_0, out8_1, out8_2, out8_3, out8_4, out8_5, out8_6, out8_7, out8_8, out8_9,
		 out9_0, out9_1, out9_2, out9_3, out9_4, out9_5, out9_6, out9_7, out9_8, out9_9,
	input [31:0]
		 W0, W1, W2, W3, W4, W5, W6, W7, W8, W9,
		 N0, N1, N2, N3, N4, N5, N6, N7, N8, N9,
	input clk, reset
);

	wire [31:0]
		ROW00__00_01, ROW00__01_02, ROW00__02_03, ROW00__03_04, ROW00__04_05, ROW00__05_06, ROW00__06_07, ROW00__07_08, ROW00__08_09, ROW00__09_10,
		ROW01__00_01, ROW01__01_02, ROW01__02_03, ROW01__03_04, ROW01__04_05, ROW01__05_06, ROW01__06_07, ROW01__07_08, ROW01__08_09, ROW01__09_10,
		ROW02__00_01, ROW02__01_02, ROW02__02_03, ROW02__03_04, ROW02__04_05, ROW02__05_06, ROW02__06_07, ROW02__07_08, ROW02__08_09, ROW02__09_10,
		ROW03__00_01, ROW03__01_02, ROW03__02_03, ROW03__03_04, ROW03__04_05, ROW03__05_06, ROW03__06_07, ROW03__07_08, ROW03__08_09, ROW03__09_10,
		ROW04__00_01, ROW04__01_02, ROW04__02_03, ROW04__03_04, ROW04__04_05, ROW04__05_06, ROW04__06_07, ROW04__07_08, ROW04__08_09, ROW04__09_10,
		ROW05__00_01, ROW05__01_02, ROW05__02_03, ROW05__03_04, ROW05__04_05, ROW05__05_06, ROW05__06_07, ROW05__07_08, ROW05__08_09, ROW05__09_10,
		ROW06__00_01, ROW06__01_02, ROW06__02_03, ROW06__03_04, ROW06__04_05, ROW06__05_06, ROW06__06_07, ROW06__07_08, ROW06__08_09, ROW06__09_10,
		ROW07__00_01, ROW07__01_02, ROW07__02_03, ROW07__03_04, ROW07__04_05, ROW07__05_06, ROW07__06_07, ROW07__07_08, ROW07__08_09, ROW07__09_10,
		ROW08__00_01, ROW08__01_02, ROW08__02_03, ROW08__03_04, ROW08__04_05, ROW08__05_06, ROW08__06_07, ROW08__07_08, ROW08__08_09, ROW08__09_10,
		ROW09__00_01, ROW09__01_02, ROW09__02_03, ROW09__03_04, ROW09__04_05, ROW09__05_06, ROW09__06_07, ROW09__07_08, ROW09__08_09, ROW09__09_10;

	wire [31:0]
		COL00__00_01, COL00__01_02, COL00__02_03, COL00__03_04, COL00__04_05, COL00__05_06, COL00__06_07, COL00__07_08, COL00__08_09, COL00__09_10,
		COL01__00_01, COL01__01_02, COL01__02_03, COL01__03_04, COL01__04_05, COL01__05_06, COL01__06_07, COL01__07_08, COL01__08_09, COL01__09_10,
		COL02__00_01, COL02__01_02, COL02__02_03, COL02__03_04, COL02__04_05, COL02__05_06, COL02__06_07, COL02__07_08, COL02__08_09, COL02__09_10,
		COL03__00_01, COL03__01_02, COL03__02_03, COL03__03_04, COL03__04_05, COL03__05_06, COL03__06_07, COL03__07_08, COL03__08_09, COL03__09_10,
		COL04__00_01, COL04__01_02, COL04__02_03, COL04__03_04, COL04__04_05, COL04__05_06, COL04__06_07, COL04__07_08, COL04__08_09, COL04__09_10,
		COL05__00_01, COL05__01_02, COL05__02_03, COL05__03_04, COL05__04_05, COL05__05_06, COL05__06_07, COL05__07_08, COL05__08_09, COL05__09_10,
		COL06__00_01, COL06__01_02, COL06__02_03, COL06__03_04, COL06__04_05, COL06__05_06, COL06__06_07, COL06__07_08, COL06__08_09, COL06__09_10,
		COL07__00_01, COL07__01_02, COL07__02_03, COL07__03_04, COL07__04_05, COL07__05_06, COL07__06_07, COL07__07_08, COL07__08_09, COL07__09_10,
		COL08__00_01, COL08__01_02, COL08__02_03, COL08__03_04, COL08__04_05, COL08__05_06, COL08__06_07, COL08__07_08, COL08__08_09, COL08__09_10,
		COL09__00_01, COL09__01_02, COL09__02_03, COL09__03_04, COL09__04_05, COL09__05_06, COL09__06_07, COL09__07_08, COL09__08_09, COL09__09_10;

	P_Element PE_00_00 {
		.out(out0_0),	.out_E(ROW00__00_01),	.out_S(COL00__00_01),
		.in_W(W0),	.in_N(N0),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_00_01 {
		.out(out0_1),	.out_E(ROW00__01_02),	.out_S(COL01__00_01),
		.in_W(W1),	.in_N(COL01__00_01),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_00_02 {
		.out(out0_2),	.out_E(ROW00__02_03),	.out_S(COL02__00_01),
		.in_W(W2),	.in_N(COL02__00_01),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_00_03 {
		.out(out0_3),	.out_E(ROW00__03_04),	.out_S(COL03__00_01),
		.in_W(W3),	.in_N(COL03__00_01),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_00_04 {
		.out(out0_4),	.out_E(ROW00__04_05),	.out_S(COL04__00_01),
		.in_W(W4),	.in_N(COL04__00_01),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_00_05 {
		.out(out0_5),	.out_E(ROW00__05_06),	.out_S(COL05__00_01),
		.in_W(W5),	.in_N(COL05__00_01),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_00_06 {
		.out(out0_6),	.out_E(ROW00__06_07),	.out_S(COL06__00_01),
		.in_W(W6),	.in_N(COL06__00_01),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_00_07 {
		.out(out0_7),	.out_E(ROW00__07_08),	.out_S(COL07__00_01),
		.in_W(W7),	.in_N(COL07__00_01),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_00_08 {
		.out(out0_8),	.out_E(ROW00__08_09),	.out_S(COL08__00_01),
		.in_W(W8),	.in_N(COL08__00_01),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_00_09 {
		.out(out0_9),	.out_E(ROW00__09_10),	.out_S(COL09__00_01),
		.in_W(W9),	.in_N(COL09__00_01),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_01_00 {
		.out(out1_0),	.out_E(ROW01__00_01),	.out_S(COL00__01_02),
		.in_W(ROW01__00_01),	.in_N(N1),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_01_01 {
		.out(out1_1),	.out_E(ROW01__01_02),	.out_S(COL01__01_02),
		.in_W(ROW01__01_02),	.in_N(COL01__01_02),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_01_02 {
		.out(out1_2),	.out_E(ROW01__02_03),	.out_S(COL02__01_02),
		.in_W(ROW01__02_03),	.in_N(COL02__01_02),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_01_03 {
		.out(out1_3),	.out_E(ROW01__03_04),	.out_S(COL03__01_02),
		.in_W(ROW01__03_04),	.in_N(COL03__01_02),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_01_04 {
		.out(out1_4),	.out_E(ROW01__04_05),	.out_S(COL04__01_02),
		.in_W(ROW01__04_05),	.in_N(COL04__01_02),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_01_05 {
		.out(out1_5),	.out_E(ROW01__05_06),	.out_S(COL05__01_02),
		.in_W(ROW01__05_06),	.in_N(COL05__01_02),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_01_06 {
		.out(out1_6),	.out_E(ROW01__06_07),	.out_S(COL06__01_02),
		.in_W(ROW01__06_07),	.in_N(COL06__01_02),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_01_07 {
		.out(out1_7),	.out_E(ROW01__07_08),	.out_S(COL07__01_02),
		.in_W(ROW01__07_08),	.in_N(COL07__01_02),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_01_08 {
		.out(out1_8),	.out_E(ROW01__08_09),	.out_S(COL08__01_02),
		.in_W(ROW01__08_09),	.in_N(COL08__01_02),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_01_09 {
		.out(out1_9),	.out_E(ROW01__09_10),	.out_S(COL09__01_02),
		.in_W(ROW01__09_10),	.in_N(COL09__01_02),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_02_00 {
		.out(out2_0),	.out_E(ROW02__00_01),	.out_S(COL00__02_03),
		.in_W(ROW02__00_01),	.in_N(N2),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_02_01 {
		.out(out2_1),	.out_E(ROW02__01_02),	.out_S(COL01__02_03),
		.in_W(ROW02__01_02),	.in_N(COL01__02_03),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_02_02 {
		.out(out2_2),	.out_E(ROW02__02_03),	.out_S(COL02__02_03),
		.in_W(ROW02__02_03),	.in_N(COL02__02_03),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_02_03 {
		.out(out2_3),	.out_E(ROW02__03_04),	.out_S(COL03__02_03),
		.in_W(ROW02__03_04),	.in_N(COL03__02_03),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_02_04 {
		.out(out2_4),	.out_E(ROW02__04_05),	.out_S(COL04__02_03),
		.in_W(ROW02__04_05),	.in_N(COL04__02_03),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_02_05 {
		.out(out2_5),	.out_E(ROW02__05_06),	.out_S(COL05__02_03),
		.in_W(ROW02__05_06),	.in_N(COL05__02_03),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_02_06 {
		.out(out2_6),	.out_E(ROW02__06_07),	.out_S(COL06__02_03),
		.in_W(ROW02__06_07),	.in_N(COL06__02_03),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_02_07 {
		.out(out2_7),	.out_E(ROW02__07_08),	.out_S(COL07__02_03),
		.in_W(ROW02__07_08),	.in_N(COL07__02_03),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_02_08 {
		.out(out2_8),	.out_E(ROW02__08_09),	.out_S(COL08__02_03),
		.in_W(ROW02__08_09),	.in_N(COL08__02_03),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_02_09 {
		.out(out2_9),	.out_E(ROW02__09_10),	.out_S(COL09__02_03),
		.in_W(ROW02__09_10),	.in_N(COL09__02_03),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_03_00 {
		.out(out3_0),	.out_E(ROW03__00_01),	.out_S(COL00__03_04),
		.in_W(ROW03__00_01),	.in_N(N3),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_03_01 {
		.out(out3_1),	.out_E(ROW03__01_02),	.out_S(COL01__03_04),
		.in_W(ROW03__01_02),	.in_N(COL01__03_04),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_03_02 {
		.out(out3_2),	.out_E(ROW03__02_03),	.out_S(COL02__03_04),
		.in_W(ROW03__02_03),	.in_N(COL02__03_04),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_03_03 {
		.out(out3_3),	.out_E(ROW03__03_04),	.out_S(COL03__03_04),
		.in_W(ROW03__03_04),	.in_N(COL03__03_04),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_03_04 {
		.out(out3_4),	.out_E(ROW03__04_05),	.out_S(COL04__03_04),
		.in_W(ROW03__04_05),	.in_N(COL04__03_04),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_03_05 {
		.out(out3_5),	.out_E(ROW03__05_06),	.out_S(COL05__03_04),
		.in_W(ROW03__05_06),	.in_N(COL05__03_04),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_03_06 {
		.out(out3_6),	.out_E(ROW03__06_07),	.out_S(COL06__03_04),
		.in_W(ROW03__06_07),	.in_N(COL06__03_04),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_03_07 {
		.out(out3_7),	.out_E(ROW03__07_08),	.out_S(COL07__03_04),
		.in_W(ROW03__07_08),	.in_N(COL07__03_04),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_03_08 {
		.out(out3_8),	.out_E(ROW03__08_09),	.out_S(COL08__03_04),
		.in_W(ROW03__08_09),	.in_N(COL08__03_04),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_03_09 {
		.out(out3_9),	.out_E(ROW03__09_10),	.out_S(COL09__03_04),
		.in_W(ROW03__09_10),	.in_N(COL09__03_04),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_04_00 {
		.out(out4_0),	.out_E(ROW04__00_01),	.out_S(COL00__04_05),
		.in_W(ROW04__00_01),	.in_N(N4),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_04_01 {
		.out(out4_1),	.out_E(ROW04__01_02),	.out_S(COL01__04_05),
		.in_W(ROW04__01_02),	.in_N(COL01__04_05),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_04_02 {
		.out(out4_2),	.out_E(ROW04__02_03),	.out_S(COL02__04_05),
		.in_W(ROW04__02_03),	.in_N(COL02__04_05),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_04_03 {
		.out(out4_3),	.out_E(ROW04__03_04),	.out_S(COL03__04_05),
		.in_W(ROW04__03_04),	.in_N(COL03__04_05),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_04_04 {
		.out(out4_4),	.out_E(ROW04__04_05),	.out_S(COL04__04_05),
		.in_W(ROW04__04_05),	.in_N(COL04__04_05),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_04_05 {
		.out(out4_5),	.out_E(ROW04__05_06),	.out_S(COL05__04_05),
		.in_W(ROW04__05_06),	.in_N(COL05__04_05),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_04_06 {
		.out(out4_6),	.out_E(ROW04__06_07),	.out_S(COL06__04_05),
		.in_W(ROW04__06_07),	.in_N(COL06__04_05),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_04_07 {
		.out(out4_7),	.out_E(ROW04__07_08),	.out_S(COL07__04_05),
		.in_W(ROW04__07_08),	.in_N(COL07__04_05),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_04_08 {
		.out(out4_8),	.out_E(ROW04__08_09),	.out_S(COL08__04_05),
		.in_W(ROW04__08_09),	.in_N(COL08__04_05),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_04_09 {
		.out(out4_9),	.out_E(ROW04__09_10),	.out_S(COL09__04_05),
		.in_W(ROW04__09_10),	.in_N(COL09__04_05),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_05_00 {
		.out(out5_0),	.out_E(ROW05__00_01),	.out_S(COL00__05_06),
		.in_W(ROW05__00_01),	.in_N(N5),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_05_01 {
		.out(out5_1),	.out_E(ROW05__01_02),	.out_S(COL01__05_06),
		.in_W(ROW05__01_02),	.in_N(COL01__05_06),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_05_02 {
		.out(out5_2),	.out_E(ROW05__02_03),	.out_S(COL02__05_06),
		.in_W(ROW05__02_03),	.in_N(COL02__05_06),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_05_03 {
		.out(out5_3),	.out_E(ROW05__03_04),	.out_S(COL03__05_06),
		.in_W(ROW05__03_04),	.in_N(COL03__05_06),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_05_04 {
		.out(out5_4),	.out_E(ROW05__04_05),	.out_S(COL04__05_06),
		.in_W(ROW05__04_05),	.in_N(COL04__05_06),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_05_05 {
		.out(out5_5),	.out_E(ROW05__05_06),	.out_S(COL05__05_06),
		.in_W(ROW05__05_06),	.in_N(COL05__05_06),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_05_06 {
		.out(out5_6),	.out_E(ROW05__06_07),	.out_S(COL06__05_06),
		.in_W(ROW05__06_07),	.in_N(COL06__05_06),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_05_07 {
		.out(out5_7),	.out_E(ROW05__07_08),	.out_S(COL07__05_06),
		.in_W(ROW05__07_08),	.in_N(COL07__05_06),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_05_08 {
		.out(out5_8),	.out_E(ROW05__08_09),	.out_S(COL08__05_06),
		.in_W(ROW05__08_09),	.in_N(COL08__05_06),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_05_09 {
		.out(out5_9),	.out_E(ROW05__09_10),	.out_S(COL09__05_06),
		.in_W(ROW05__09_10),	.in_N(COL09__05_06),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_06_00 {
		.out(out6_0),	.out_E(ROW06__00_01),	.out_S(COL00__06_07),
		.in_W(ROW06__00_01),	.in_N(N6),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_06_01 {
		.out(out6_1),	.out_E(ROW06__01_02),	.out_S(COL01__06_07),
		.in_W(ROW06__01_02),	.in_N(COL01__06_07),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_06_02 {
		.out(out6_2),	.out_E(ROW06__02_03),	.out_S(COL02__06_07),
		.in_W(ROW06__02_03),	.in_N(COL02__06_07),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_06_03 {
		.out(out6_3),	.out_E(ROW06__03_04),	.out_S(COL03__06_07),
		.in_W(ROW06__03_04),	.in_N(COL03__06_07),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_06_04 {
		.out(out6_4),	.out_E(ROW06__04_05),	.out_S(COL04__06_07),
		.in_W(ROW06__04_05),	.in_N(COL04__06_07),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_06_05 {
		.out(out6_5),	.out_E(ROW06__05_06),	.out_S(COL05__06_07),
		.in_W(ROW06__05_06),	.in_N(COL05__06_07),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_06_06 {
		.out(out6_6),	.out_E(ROW06__06_07),	.out_S(COL06__06_07),
		.in_W(ROW06__06_07),	.in_N(COL06__06_07),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_06_07 {
		.out(out6_7),	.out_E(ROW06__07_08),	.out_S(COL07__06_07),
		.in_W(ROW06__07_08),	.in_N(COL07__06_07),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_06_08 {
		.out(out6_8),	.out_E(ROW06__08_09),	.out_S(COL08__06_07),
		.in_W(ROW06__08_09),	.in_N(COL08__06_07),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_06_09 {
		.out(out6_9),	.out_E(ROW06__09_10),	.out_S(COL09__06_07),
		.in_W(ROW06__09_10),	.in_N(COL09__06_07),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_07_00 {
		.out(out7_0),	.out_E(ROW07__00_01),	.out_S(COL00__07_08),
		.in_W(ROW07__00_01),	.in_N(N7),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_07_01 {
		.out(out7_1),	.out_E(ROW07__01_02),	.out_S(COL01__07_08),
		.in_W(ROW07__01_02),	.in_N(COL01__07_08),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_07_02 {
		.out(out7_2),	.out_E(ROW07__02_03),	.out_S(COL02__07_08),
		.in_W(ROW07__02_03),	.in_N(COL02__07_08),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_07_03 {
		.out(out7_3),	.out_E(ROW07__03_04),	.out_S(COL03__07_08),
		.in_W(ROW07__03_04),	.in_N(COL03__07_08),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_07_04 {
		.out(out7_4),	.out_E(ROW07__04_05),	.out_S(COL04__07_08),
		.in_W(ROW07__04_05),	.in_N(COL04__07_08),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_07_05 {
		.out(out7_5),	.out_E(ROW07__05_06),	.out_S(COL05__07_08),
		.in_W(ROW07__05_06),	.in_N(COL05__07_08),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_07_06 {
		.out(out7_6),	.out_E(ROW07__06_07),	.out_S(COL06__07_08),
		.in_W(ROW07__06_07),	.in_N(COL06__07_08),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_07_07 {
		.out(out7_7),	.out_E(ROW07__07_08),	.out_S(COL07__07_08),
		.in_W(ROW07__07_08),	.in_N(COL07__07_08),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_07_08 {
		.out(out7_8),	.out_E(ROW07__08_09),	.out_S(COL08__07_08),
		.in_W(ROW07__08_09),	.in_N(COL08__07_08),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_07_09 {
		.out(out7_9),	.out_E(ROW07__09_10),	.out_S(COL09__07_08),
		.in_W(ROW07__09_10),	.in_N(COL09__07_08),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_08_00 {
		.out(out8_0),	.out_E(ROW08__00_01),	.out_S(COL00__08_09),
		.in_W(ROW08__00_01),	.in_N(N8),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_08_01 {
		.out(out8_1),	.out_E(ROW08__01_02),	.out_S(COL01__08_09),
		.in_W(ROW08__01_02),	.in_N(COL01__08_09),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_08_02 {
		.out(out8_2),	.out_E(ROW08__02_03),	.out_S(COL02__08_09),
		.in_W(ROW08__02_03),	.in_N(COL02__08_09),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_08_03 {
		.out(out8_3),	.out_E(ROW08__03_04),	.out_S(COL03__08_09),
		.in_W(ROW08__03_04),	.in_N(COL03__08_09),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_08_04 {
		.out(out8_4),	.out_E(ROW08__04_05),	.out_S(COL04__08_09),
		.in_W(ROW08__04_05),	.in_N(COL04__08_09),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_08_05 {
		.out(out8_5),	.out_E(ROW08__05_06),	.out_S(COL05__08_09),
		.in_W(ROW08__05_06),	.in_N(COL05__08_09),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_08_06 {
		.out(out8_6),	.out_E(ROW08__06_07),	.out_S(COL06__08_09),
		.in_W(ROW08__06_07),	.in_N(COL06__08_09),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_08_07 {
		.out(out8_7),	.out_E(ROW08__07_08),	.out_S(COL07__08_09),
		.in_W(ROW08__07_08),	.in_N(COL07__08_09),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_08_08 {
		.out(out8_8),	.out_E(ROW08__08_09),	.out_S(COL08__08_09),
		.in_W(ROW08__08_09),	.in_N(COL08__08_09),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_08_09 {
		.out(out8_9),	.out_E(ROW08__09_10),	.out_S(COL09__08_09),
		.in_W(ROW08__09_10),	.in_N(COL09__08_09),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_09_00 {
		.out(out9_0),	.out_E(ROW09__00_01),	.out_S(COL00__09_10),
		.in_W(ROW09__00_01),	.in_N(N9),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_09_01 {
		.out(out9_1),	.out_E(ROW09__01_02),	.out_S(COL01__09_10),
		.in_W(ROW09__01_02),	.in_N(COL01__09_10),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_09_02 {
		.out(out9_2),	.out_E(ROW09__02_03),	.out_S(COL02__09_10),
		.in_W(ROW09__02_03),	.in_N(COL02__09_10),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_09_03 {
		.out(out9_3),	.out_E(ROW09__03_04),	.out_S(COL03__09_10),
		.in_W(ROW09__03_04),	.in_N(COL03__09_10),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_09_04 {
		.out(out9_4),	.out_E(ROW09__04_05),	.out_S(COL04__09_10),
		.in_W(ROW09__04_05),	.in_N(COL04__09_10),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_09_05 {
		.out(out9_5),	.out_E(ROW09__05_06),	.out_S(COL05__09_10),
		.in_W(ROW09__05_06),	.in_N(COL05__09_10),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_09_06 {
		.out(out9_6),	.out_E(ROW09__06_07),	.out_S(COL06__09_10),
		.in_W(ROW09__06_07),	.in_N(COL06__09_10),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_09_07 {
		.out(out9_7),	.out_E(ROW09__07_08),	.out_S(COL07__09_10),
		.in_W(ROW09__07_08),	.in_N(COL07__09_10),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_09_08 {
		.out(out9_8),	.out_E(ROW09__08_09),	.out_S(COL08__09_10),
		.in_W(ROW09__08_09),	.in_N(COL08__09_10),
		.clk(clk),	.reset(reset)
	};
	P_Element PE_09_09 {
		.out(out9_9),	.out_E(ROW09__09_10),	.out_S(COL09__09_10),
		.in_W(ROW09__09_10),	.in_N(COL09__09_10),
		.clk(clk),	.reset(reset)
	};
endmodule
