module Systolic_Array10x10 (
	output [31:0]
		 out0_0, out0_1, out0_2, out0_3, out0_4, out0_5, out0_6, out0_7, out0_8, out0_9,
		 out1_0, out1_1, out1_2, out1_3, out1_4, out1_5, out1_6, out1_7, out1_8, out1_9,
		 out2_0, out2_1, out2_2, out2_3, out2_4, out2_5, out2_6, out2_7, out2_8, out2_9,
		 out3_0, out3_1, out3_2, out3_3, out3_4, out3_5, out3_6, out3_7, out3_8, out3_9,
		 out4_0, out4_1, out4_2, out4_3, out4_4, out4_5, out4_6, out4_7, out4_8, out4_9,
		 out5_0, out5_1, out5_2, out5_3, out5_4, out5_5, out5_6, out5_7, out5_8, out5_9,
		 out6_0, out6_1, out6_2, out6_3, out6_4, out6_5, out6_6, out6_7, out6_8, out6_9,
		 out7_0, out7_1, out7_2, out7_3, out7_4, out7_5, out7_6, out7_7, out7_8, out7_9,
		 out8_0, out8_1, out8_2, out8_3, out8_4, out8_5, out8_6, out8_7, out8_8, out8_9,
		 out9_0, out9_1, out9_2, out9_3, out9_4, out9_5, out9_6, out9_7, out9_8, out9_9,
	input [31:0]
		 W0, W1, W2, W3, W4, W5, W6, W7, W8, W9,
		 N0, N1, N2, N3, N4, N5, N6, N7, N8, N9,
	input clk, reset
);

	wire [31:0]
		ROW00_00, ROW00_01, ROW00_02, ROW00_03, ROW00_04, ROW00_05, ROW00_06, ROW00_07, ROW00_08, ROW00_09,
		ROW01_00, ROW01_01, ROW01_02, ROW01_03, ROW01_04, ROW01_05, ROW01_06, ROW01_07, ROW01_08, ROW01_09,
		ROW02_00, ROW02_01, ROW02_02, ROW02_03, ROW02_04, ROW02_05, ROW02_06, ROW02_07, ROW02_08, ROW02_09,
		ROW03_00, ROW03_01, ROW03_02, ROW03_03, ROW03_04, ROW03_05, ROW03_06, ROW03_07, ROW03_08, ROW03_09,
		ROW04_00, ROW04_01, ROW04_02, ROW04_03, ROW04_04, ROW04_05, ROW04_06, ROW04_07, ROW04_08, ROW04_09,
		ROW05_00, ROW05_01, ROW05_02, ROW05_03, ROW05_04, ROW05_05, ROW05_06, ROW05_07, ROW05_08, ROW05_09,
		ROW06_00, ROW06_01, ROW06_02, ROW06_03, ROW06_04, ROW06_05, ROW06_06, ROW06_07, ROW06_08, ROW06_09,
		ROW07_00, ROW07_01, ROW07_02, ROW07_03, ROW07_04, ROW07_05, ROW07_06, ROW07_07, ROW07_08, ROW07_09,
		ROW08_00, ROW08_01, ROW08_02, ROW08_03, ROW08_04, ROW08_05, ROW08_06, ROW08_07, ROW08_08, ROW08_09,
		ROW09_00, ROW09_01, ROW09_02, ROW09_03, ROW09_04, ROW09_05, ROW09_06, ROW09_07, ROW09_08, ROW09_09;

	wire [31:0]
		COL00_00, COL00_01, COL00_02, COL00_03, COL00_04, COL00_05, COL00_06, COL00_07, COL00_08, COL00_09,
		COL01_00, COL01_01, COL01_02, COL01_03, COL01_04, COL01_05, COL01_06, COL01_07, COL01_08, COL01_09,
		COL02_00, COL02_01, COL02_02, COL02_03, COL02_04, COL02_05, COL02_06, COL02_07, COL02_08, COL02_09,
		COL03_00, COL03_01, COL03_02, COL03_03, COL03_04, COL03_05, COL03_06, COL03_07, COL03_08, COL03_09,
		COL04_00, COL04_01, COL04_02, COL04_03, COL04_04, COL04_05, COL04_06, COL04_07, COL04_08, COL04_09,
		COL05_00, COL05_01, COL05_02, COL05_03, COL05_04, COL05_05, COL05_06, COL05_07, COL05_08, COL05_09,
		COL06_00, COL06_01, COL06_02, COL06_03, COL06_04, COL06_05, COL06_06, COL06_07, COL06_08, COL06_09,
		COL07_00, COL07_01, COL07_02, COL07_03, COL07_04, COL07_05, COL07_06, COL07_07, COL07_08, COL07_09,
		COL08_00, COL08_01, COL08_02, COL08_03, COL08_04, COL08_05, COL08_06, COL08_07, COL08_08, COL08_09,
		COL09_00, COL09_01, COL09_02, COL09_03, COL09_04, COL09_05, COL09_06, COL09_07, COL09_08, COL09_09;

	P_Element PE_00_00 (
		.OUT(out0_0),	.OUT_RIGHT(ROW00_00),	.OUT_BOTTOM(COL00_00),
		.IN_LEFT(W0),	.IN_TOP(N0),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_00_01 (
		.OUT(out0_1),	.OUT_RIGHT(ROW00_01),	.OUT_BOTTOM(COL00_01),
		.IN_LEFT(ROW00_00),	.IN_TOP(N1),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_00_02 (
		.OUT(out0_2),	.OUT_RIGHT(ROW00_02),	.OUT_BOTTOM(COL00_02),
		.IN_LEFT(ROW00_01),	.IN_TOP(N2),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_00_03 (
		.OUT(out0_3),	.OUT_RIGHT(ROW00_03),	.OUT_BOTTOM(COL00_03),
		.IN_LEFT(ROW00_02),	.IN_TOP(N3),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_00_04 (
		.OUT(out0_4),	.OUT_RIGHT(ROW00_04),	.OUT_BOTTOM(COL00_04),
		.IN_LEFT(ROW00_03),	.IN_TOP(N4),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_00_05 (
		.OUT(out0_5),	.OUT_RIGHT(ROW00_05),	.OUT_BOTTOM(COL00_05),
		.IN_LEFT(ROW00_04),	.IN_TOP(N5),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_00_06 (
		.OUT(out0_6),	.OUT_RIGHT(ROW00_06),	.OUT_BOTTOM(COL00_06),
		.IN_LEFT(ROW00_05),	.IN_TOP(N6),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_00_07 (
		.OUT(out0_7),	.OUT_RIGHT(ROW00_07),	.OUT_BOTTOM(COL00_07),
		.IN_LEFT(ROW00_06),	.IN_TOP(N7),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_00_08 (
		.OUT(out0_8),	.OUT_RIGHT(ROW00_08),	.OUT_BOTTOM(COL00_08),
		.IN_LEFT(ROW00_07),	.IN_TOP(N8),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_00_09 (
		.OUT(out0_9),	.OUT_RIGHT(ROW00_09),	.OUT_BOTTOM(COL00_09),
		.IN_LEFT(ROW00_08),	.IN_TOP(N9),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_01_00 (
		.OUT(out1_0),	.OUT_RIGHT(ROW01_00),	.OUT_BOTTOM(COL01_00),
		.IN_LEFT(W1),	.IN_TOP(COL00_00),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_01_01 (
		.OUT(out1_1),	.OUT_RIGHT(ROW01_01),	.OUT_BOTTOM(COL01_01),
		.IN_LEFT(ROW01_00),	.IN_TOP(COL00_01),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_01_02 (
		.OUT(out1_2),	.OUT_RIGHT(ROW01_02),	.OUT_BOTTOM(COL01_02),
		.IN_LEFT(ROW01_01),	.IN_TOP(COL00_02),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_01_03 (
		.OUT(out1_3),	.OUT_RIGHT(ROW01_03),	.OUT_BOTTOM(COL01_03),
		.IN_LEFT(ROW01_02),	.IN_TOP(COL00_03),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_01_04 (
		.OUT(out1_4),	.OUT_RIGHT(ROW01_04),	.OUT_BOTTOM(COL01_04),
		.IN_LEFT(ROW01_03),	.IN_TOP(COL00_04),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_01_05 (
		.OUT(out1_5),	.OUT_RIGHT(ROW01_05),	.OUT_BOTTOM(COL01_05),
		.IN_LEFT(ROW01_04),	.IN_TOP(COL00_05),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_01_06 (
		.OUT(out1_6),	.OUT_RIGHT(ROW01_06),	.OUT_BOTTOM(COL01_06),
		.IN_LEFT(ROW01_05),	.IN_TOP(COL00_06),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_01_07 (
		.OUT(out1_7),	.OUT_RIGHT(ROW01_07),	.OUT_BOTTOM(COL01_07),
		.IN_LEFT(ROW01_06),	.IN_TOP(COL00_07),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_01_08 (
		.OUT(out1_8),	.OUT_RIGHT(ROW01_08),	.OUT_BOTTOM(COL01_08),
		.IN_LEFT(ROW01_07),	.IN_TOP(COL00_08),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_01_09 (
		.OUT(out1_9),	.OUT_RIGHT(ROW01_09),	.OUT_BOTTOM(COL01_09),
		.IN_LEFT(ROW01_08),	.IN_TOP(COL00_09),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_02_00 (
		.OUT(out2_0),	.OUT_RIGHT(ROW02_00),	.OUT_BOTTOM(COL02_00),
		.IN_LEFT(W2),	.IN_TOP(COL01_00),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_02_01 (
		.OUT(out2_1),	.OUT_RIGHT(ROW02_01),	.OUT_BOTTOM(COL02_01),
		.IN_LEFT(ROW02_00),	.IN_TOP(COL01_01),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_02_02 (
		.OUT(out2_2),	.OUT_RIGHT(ROW02_02),	.OUT_BOTTOM(COL02_02),
		.IN_LEFT(ROW02_01),	.IN_TOP(COL01_02),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_02_03 (
		.OUT(out2_3),	.OUT_RIGHT(ROW02_03),	.OUT_BOTTOM(COL02_03),
		.IN_LEFT(ROW02_02),	.IN_TOP(COL01_03),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_02_04 (
		.OUT(out2_4),	.OUT_RIGHT(ROW02_04),	.OUT_BOTTOM(COL02_04),
		.IN_LEFT(ROW02_03),	.IN_TOP(COL01_04),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_02_05 (
		.OUT(out2_5),	.OUT_RIGHT(ROW02_05),	.OUT_BOTTOM(COL02_05),
		.IN_LEFT(ROW02_04),	.IN_TOP(COL01_05),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_02_06 (
		.OUT(out2_6),	.OUT_RIGHT(ROW02_06),	.OUT_BOTTOM(COL02_06),
		.IN_LEFT(ROW02_05),	.IN_TOP(COL01_06),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_02_07 (
		.OUT(out2_7),	.OUT_RIGHT(ROW02_07),	.OUT_BOTTOM(COL02_07),
		.IN_LEFT(ROW02_06),	.IN_TOP(COL01_07),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_02_08 (
		.OUT(out2_8),	.OUT_RIGHT(ROW02_08),	.OUT_BOTTOM(COL02_08),
		.IN_LEFT(ROW02_07),	.IN_TOP(COL01_08),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_02_09 (
		.OUT(out2_9),	.OUT_RIGHT(ROW02_09),	.OUT_BOTTOM(COL02_09),
		.IN_LEFT(ROW02_08),	.IN_TOP(COL01_09),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_03_00 (
		.OUT(out3_0),	.OUT_RIGHT(ROW03_00),	.OUT_BOTTOM(COL03_00),
		.IN_LEFT(W3),	.IN_TOP(COL02_00),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_03_01 (
		.OUT(out3_1),	.OUT_RIGHT(ROW03_01),	.OUT_BOTTOM(COL03_01),
		.IN_LEFT(ROW03_00),	.IN_TOP(COL02_01),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_03_02 (
		.OUT(out3_2),	.OUT_RIGHT(ROW03_02),	.OUT_BOTTOM(COL03_02),
		.IN_LEFT(ROW03_01),	.IN_TOP(COL02_02),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_03_03 (
		.OUT(out3_3),	.OUT_RIGHT(ROW03_03),	.OUT_BOTTOM(COL03_03),
		.IN_LEFT(ROW03_02),	.IN_TOP(COL02_03),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_03_04 (
		.OUT(out3_4),	.OUT_RIGHT(ROW03_04),	.OUT_BOTTOM(COL03_04),
		.IN_LEFT(ROW03_03),	.IN_TOP(COL02_04),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_03_05 (
		.OUT(out3_5),	.OUT_RIGHT(ROW03_05),	.OUT_BOTTOM(COL03_05),
		.IN_LEFT(ROW03_04),	.IN_TOP(COL02_05),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_03_06 (
		.OUT(out3_6),	.OUT_RIGHT(ROW03_06),	.OUT_BOTTOM(COL03_06),
		.IN_LEFT(ROW03_05),	.IN_TOP(COL02_06),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_03_07 (
		.OUT(out3_7),	.OUT_RIGHT(ROW03_07),	.OUT_BOTTOM(COL03_07),
		.IN_LEFT(ROW03_06),	.IN_TOP(COL02_07),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_03_08 (
		.OUT(out3_8),	.OUT_RIGHT(ROW03_08),	.OUT_BOTTOM(COL03_08),
		.IN_LEFT(ROW03_07),	.IN_TOP(COL02_08),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_03_09 (
		.OUT(out3_9),	.OUT_RIGHT(ROW03_09),	.OUT_BOTTOM(COL03_09),
		.IN_LEFT(ROW03_08),	.IN_TOP(COL02_09),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_04_00 (
		.OUT(out4_0),	.OUT_RIGHT(ROW04_00),	.OUT_BOTTOM(COL04_00),
		.IN_LEFT(W4),	.IN_TOP(COL03_00),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_04_01 (
		.OUT(out4_1),	.OUT_RIGHT(ROW04_01),	.OUT_BOTTOM(COL04_01),
		.IN_LEFT(ROW04_00),	.IN_TOP(COL03_01),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_04_02 (
		.OUT(out4_2),	.OUT_RIGHT(ROW04_02),	.OUT_BOTTOM(COL04_02),
		.IN_LEFT(ROW04_01),	.IN_TOP(COL03_02),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_04_03 (
		.OUT(out4_3),	.OUT_RIGHT(ROW04_03),	.OUT_BOTTOM(COL04_03),
		.IN_LEFT(ROW04_02),	.IN_TOP(COL03_03),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_04_04 (
		.OUT(out4_4),	.OUT_RIGHT(ROW04_04),	.OUT_BOTTOM(COL04_04),
		.IN_LEFT(ROW04_03),	.IN_TOP(COL03_04),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_04_05 (
		.OUT(out4_5),	.OUT_RIGHT(ROW04_05),	.OUT_BOTTOM(COL04_05),
		.IN_LEFT(ROW04_04),	.IN_TOP(COL03_05),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_04_06 (
		.OUT(out4_6),	.OUT_RIGHT(ROW04_06),	.OUT_BOTTOM(COL04_06),
		.IN_LEFT(ROW04_05),	.IN_TOP(COL03_06),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_04_07 (
		.OUT(out4_7),	.OUT_RIGHT(ROW04_07),	.OUT_BOTTOM(COL04_07),
		.IN_LEFT(ROW04_06),	.IN_TOP(COL03_07),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_04_08 (
		.OUT(out4_8),	.OUT_RIGHT(ROW04_08),	.OUT_BOTTOM(COL04_08),
		.IN_LEFT(ROW04_07),	.IN_TOP(COL03_08),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_04_09 (
		.OUT(out4_9),	.OUT_RIGHT(ROW04_09),	.OUT_BOTTOM(COL04_09),
		.IN_LEFT(ROW04_08),	.IN_TOP(COL03_09),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_05_00 (
		.OUT(out5_0),	.OUT_RIGHT(ROW05_00),	.OUT_BOTTOM(COL05_00),
		.IN_LEFT(W5),	.IN_TOP(COL04_00),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_05_01 (
		.OUT(out5_1),	.OUT_RIGHT(ROW05_01),	.OUT_BOTTOM(COL05_01),
		.IN_LEFT(ROW05_00),	.IN_TOP(COL04_01),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_05_02 (
		.OUT(out5_2),	.OUT_RIGHT(ROW05_02),	.OUT_BOTTOM(COL05_02),
		.IN_LEFT(ROW05_01),	.IN_TOP(COL04_02),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_05_03 (
		.OUT(out5_3),	.OUT_RIGHT(ROW05_03),	.OUT_BOTTOM(COL05_03),
		.IN_LEFT(ROW05_02),	.IN_TOP(COL04_03),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_05_04 (
		.OUT(out5_4),	.OUT_RIGHT(ROW05_04),	.OUT_BOTTOM(COL05_04),
		.IN_LEFT(ROW05_03),	.IN_TOP(COL04_04),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_05_05 (
		.OUT(out5_5),	.OUT_RIGHT(ROW05_05),	.OUT_BOTTOM(COL05_05),
		.IN_LEFT(ROW05_04),	.IN_TOP(COL04_05),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_05_06 (
		.OUT(out5_6),	.OUT_RIGHT(ROW05_06),	.OUT_BOTTOM(COL05_06),
		.IN_LEFT(ROW05_05),	.IN_TOP(COL04_06),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_05_07 (
		.OUT(out5_7),	.OUT_RIGHT(ROW05_07),	.OUT_BOTTOM(COL05_07),
		.IN_LEFT(ROW05_06),	.IN_TOP(COL04_07),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_05_08 (
		.OUT(out5_8),	.OUT_RIGHT(ROW05_08),	.OUT_BOTTOM(COL05_08),
		.IN_LEFT(ROW05_07),	.IN_TOP(COL04_08),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_05_09 (
		.OUT(out5_9),	.OUT_RIGHT(ROW05_09),	.OUT_BOTTOM(COL05_09),
		.IN_LEFT(ROW05_08),	.IN_TOP(COL04_09),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_06_00 (
		.OUT(out6_0),	.OUT_RIGHT(ROW06_00),	.OUT_BOTTOM(COL06_00),
		.IN_LEFT(W6),	.IN_TOP(COL05_00),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_06_01 (
		.OUT(out6_1),	.OUT_RIGHT(ROW06_01),	.OUT_BOTTOM(COL06_01),
		.IN_LEFT(ROW06_00),	.IN_TOP(COL05_01),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_06_02 (
		.OUT(out6_2),	.OUT_RIGHT(ROW06_02),	.OUT_BOTTOM(COL06_02),
		.IN_LEFT(ROW06_01),	.IN_TOP(COL05_02),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_06_03 (
		.OUT(out6_3),	.OUT_RIGHT(ROW06_03),	.OUT_BOTTOM(COL06_03),
		.IN_LEFT(ROW06_02),	.IN_TOP(COL05_03),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_06_04 (
		.OUT(out6_4),	.OUT_RIGHT(ROW06_04),	.OUT_BOTTOM(COL06_04),
		.IN_LEFT(ROW06_03),	.IN_TOP(COL05_04),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_06_05 (
		.OUT(out6_5),	.OUT_RIGHT(ROW06_05),	.OUT_BOTTOM(COL06_05),
		.IN_LEFT(ROW06_04),	.IN_TOP(COL05_05),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_06_06 (
		.OUT(out6_6),	.OUT_RIGHT(ROW06_06),	.OUT_BOTTOM(COL06_06),
		.IN_LEFT(ROW06_05),	.IN_TOP(COL05_06),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_06_07 (
		.OUT(out6_7),	.OUT_RIGHT(ROW06_07),	.OUT_BOTTOM(COL06_07),
		.IN_LEFT(ROW06_06),	.IN_TOP(COL05_07),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_06_08 (
		.OUT(out6_8),	.OUT_RIGHT(ROW06_08),	.OUT_BOTTOM(COL06_08),
		.IN_LEFT(ROW06_07),	.IN_TOP(COL05_08),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_06_09 (
		.OUT(out6_9),	.OUT_RIGHT(ROW06_09),	.OUT_BOTTOM(COL06_09),
		.IN_LEFT(ROW06_08),	.IN_TOP(COL05_09),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_07_00 (
		.OUT(out7_0),	.OUT_RIGHT(ROW07_00),	.OUT_BOTTOM(COL07_00),
		.IN_LEFT(W7),	.IN_TOP(COL06_00),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_07_01 (
		.OUT(out7_1),	.OUT_RIGHT(ROW07_01),	.OUT_BOTTOM(COL07_01),
		.IN_LEFT(ROW07_00),	.IN_TOP(COL06_01),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_07_02 (
		.OUT(out7_2),	.OUT_RIGHT(ROW07_02),	.OUT_BOTTOM(COL07_02),
		.IN_LEFT(ROW07_01),	.IN_TOP(COL06_02),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_07_03 (
		.OUT(out7_3),	.OUT_RIGHT(ROW07_03),	.OUT_BOTTOM(COL07_03),
		.IN_LEFT(ROW07_02),	.IN_TOP(COL06_03),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_07_04 (
		.OUT(out7_4),	.OUT_RIGHT(ROW07_04),	.OUT_BOTTOM(COL07_04),
		.IN_LEFT(ROW07_03),	.IN_TOP(COL06_04),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_07_05 (
		.OUT(out7_5),	.OUT_RIGHT(ROW07_05),	.OUT_BOTTOM(COL07_05),
		.IN_LEFT(ROW07_04),	.IN_TOP(COL06_05),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_07_06 (
		.OUT(out7_6),	.OUT_RIGHT(ROW07_06),	.OUT_BOTTOM(COL07_06),
		.IN_LEFT(ROW07_05),	.IN_TOP(COL06_06),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_07_07 (
		.OUT(out7_7),	.OUT_RIGHT(ROW07_07),	.OUT_BOTTOM(COL07_07),
		.IN_LEFT(ROW07_06),	.IN_TOP(COL06_07),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_07_08 (
		.OUT(out7_8),	.OUT_RIGHT(ROW07_08),	.OUT_BOTTOM(COL07_08),
		.IN_LEFT(ROW07_07),	.IN_TOP(COL06_08),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_07_09 (
		.OUT(out7_9),	.OUT_RIGHT(ROW07_09),	.OUT_BOTTOM(COL07_09),
		.IN_LEFT(ROW07_08),	.IN_TOP(COL06_09),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_08_00 (
		.OUT(out8_0),	.OUT_RIGHT(ROW08_00),	.OUT_BOTTOM(COL08_00),
		.IN_LEFT(W8),	.IN_TOP(COL07_00),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_08_01 (
		.OUT(out8_1),	.OUT_RIGHT(ROW08_01),	.OUT_BOTTOM(COL08_01),
		.IN_LEFT(ROW08_00),	.IN_TOP(COL07_01),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_08_02 (
		.OUT(out8_2),	.OUT_RIGHT(ROW08_02),	.OUT_BOTTOM(COL08_02),
		.IN_LEFT(ROW08_01),	.IN_TOP(COL07_02),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_08_03 (
		.OUT(out8_3),	.OUT_RIGHT(ROW08_03),	.OUT_BOTTOM(COL08_03),
		.IN_LEFT(ROW08_02),	.IN_TOP(COL07_03),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_08_04 (
		.OUT(out8_4),	.OUT_RIGHT(ROW08_04),	.OUT_BOTTOM(COL08_04),
		.IN_LEFT(ROW08_03),	.IN_TOP(COL07_04),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_08_05 (
		.OUT(out8_5),	.OUT_RIGHT(ROW08_05),	.OUT_BOTTOM(COL08_05),
		.IN_LEFT(ROW08_04),	.IN_TOP(COL07_05),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_08_06 (
		.OUT(out8_6),	.OUT_RIGHT(ROW08_06),	.OUT_BOTTOM(COL08_06),
		.IN_LEFT(ROW08_05),	.IN_TOP(COL07_06),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_08_07 (
		.OUT(out8_7),	.OUT_RIGHT(ROW08_07),	.OUT_BOTTOM(COL08_07),
		.IN_LEFT(ROW08_06),	.IN_TOP(COL07_07),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_08_08 (
		.OUT(out8_8),	.OUT_RIGHT(ROW08_08),	.OUT_BOTTOM(COL08_08),
		.IN_LEFT(ROW08_07),	.IN_TOP(COL07_08),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_08_09 (
		.OUT(out8_9),	.OUT_RIGHT(ROW08_09),	.OUT_BOTTOM(COL08_09),
		.IN_LEFT(ROW08_08),	.IN_TOP(COL07_09),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_09_00 (
		.OUT(out9_0),	.OUT_RIGHT(ROW09_00),	.OUT_BOTTOM(COL09_00),
		.IN_LEFT(W9),	.IN_TOP(COL08_00),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_09_01 (
		.OUT(out9_1),	.OUT_RIGHT(ROW09_01),	.OUT_BOTTOM(COL09_01),
		.IN_LEFT(ROW09_00),	.IN_TOP(COL08_01),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_09_02 (
		.OUT(out9_2),	.OUT_RIGHT(ROW09_02),	.OUT_BOTTOM(COL09_02),
		.IN_LEFT(ROW09_01),	.IN_TOP(COL08_02),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_09_03 (
		.OUT(out9_3),	.OUT_RIGHT(ROW09_03),	.OUT_BOTTOM(COL09_03),
		.IN_LEFT(ROW09_02),	.IN_TOP(COL08_03),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_09_04 (
		.OUT(out9_4),	.OUT_RIGHT(ROW09_04),	.OUT_BOTTOM(COL09_04),
		.IN_LEFT(ROW09_03),	.IN_TOP(COL08_04),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_09_05 (
		.OUT(out9_5),	.OUT_RIGHT(ROW09_05),	.OUT_BOTTOM(COL09_05),
		.IN_LEFT(ROW09_04),	.IN_TOP(COL08_05),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_09_06 (
		.OUT(out9_6),	.OUT_RIGHT(ROW09_06),	.OUT_BOTTOM(COL09_06),
		.IN_LEFT(ROW09_05),	.IN_TOP(COL08_06),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_09_07 (
		.OUT(out9_7),	.OUT_RIGHT(ROW09_07),	.OUT_BOTTOM(COL09_07),
		.IN_LEFT(ROW09_06),	.IN_TOP(COL08_07),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_09_08 (
		.OUT(out9_8),	.OUT_RIGHT(ROW09_08),	.OUT_BOTTOM(COL09_08),
		.IN_LEFT(ROW09_07),	.IN_TOP(COL08_08),
		.CLK(clk),	.RST_N(reset)
	);
	P_Element PE_09_09 (
		.OUT(out9_9),	.OUT_RIGHT(ROW09_09),	.OUT_BOTTOM(COL09_09),
		.IN_LEFT(ROW09_08),	.IN_TOP(COL08_09),
		.CLK(clk),	.RST_N(reset)
	);
endmodule
